create keyspace Indexing;

use Indexing;

create column family Configuration
  with comparator = 'UTF8Type'
  and default_validation_class = 'UTF8Type'
  and key_validation_class = 'UTF8Type';

create column family Indexes
  with comparator = 'CompositeType(UTF8Type, UTF8Type, UTF8Type, UTF8Type, UTF8Type)'
  and default_validation_class = 'UTF8Type'
  and key_validation_class = 'UTF8Type';
